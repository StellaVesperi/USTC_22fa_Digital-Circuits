module d_ff_r(  
input clk,rst_n,d,  
output reg q);  
	always@(posedge clk)  
	begin  
		if(rst_n==0)  
			q <= 1'b0;  
		else  
			q <= d;  
	end  
endmodule