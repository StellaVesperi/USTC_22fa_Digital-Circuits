module d_ff(
    input clk, d,
    output reg q);
    always @ (posedge clk)
        q <= d;
endmodule

/*˵���� reg�� always �� posedge �� Verilog �еĹؼ��֣� ���� always ��ʾ����Ǹ��������顣
reg ��ǰ��ѧϰ���� wire �ؼ������ƣ���һ���������ͣ���Ϊ�Ĵ������͡�
���ڳ�ѧ�ߣ����Լ򵥵����Ϊ������ always �����ڱ���ֵ���źţ���Ӧ����Ϊ reg ���͡� 
posedge Ϊ�¼����ƹؼ��֣� ��������еġ�posedge clk����ʾ��clk �źŵ������ء���һ�¼���
���⣬��ʱ���߼���·�У��źŸ�ֵ���á�<=������������ֵ�� ,�����ǡ�=����������ֵ���� 
�����ָ�ֵ��ʽ�������ݲ����ܣ�����ֻ���סһ��ԭ������߼�����������ֵ��=����ʱ���߼����÷�������ֵ��<=�� ��
*/
