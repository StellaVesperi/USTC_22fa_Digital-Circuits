//��ʱ���źŵ������ز������õĴ������ĸ�λ�ź�
// Called ͬ����λ
module d_ff_r_syn(
    input clk, rst_n, d,
    output reg q);
    always @ (posedge clk)
    begin
        if (rst_n == 0)
            q <= 1'b0;
        else 
            q <= d;
    end
endmodule

/*
˵������δ��������³����� begin�� end�� if�� else �ĸ��ؼ��֣�
���� begin/end����ɶԳ��֣����ڱ���������������䣬
�����������У� begin/end ֮��Ĵ��붼����ͬһ always �顣 
if�� else ���������жϣ��ںܶ����������ж��г��֣��京��Ҳ��һ�����˴�����׸���� 
��1��b0����һ�����ݱ�ʾ��ʽ��һ���ʽΪ������λ��������ֵ����
�����б�ʾ����һ�� 1bit �����ݣ��ö����Ʊ�ʾ����ֵΪ 0��
*/
